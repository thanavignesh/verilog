library verilog;
use verilog.vl_types.all;
entity srtb is
end srtb;
