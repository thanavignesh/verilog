library verilog;
use verilog.vl_types.all;
entity jktb is
end jktb;
