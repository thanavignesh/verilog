library verilog;
use verilog.vl_types.all;
entity binarytb is
end binarytb;
