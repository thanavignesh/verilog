library verilog;
use verilog.vl_types.all;
entity asynctb is
end asynctb;
