library verilog;
use verilog.vl_types.all;
entity bcdtb is
end bcdtb;
