library verilog;
use verilog.vl_types.all;
entity syntb is
end syntb;
