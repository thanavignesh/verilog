library verilog;
use verilog.vl_types.all;
entity tff_tb is
end tff_tb;
